`define WORD_SIZE 16 
`define ADDR_SIZE 8
