`define WORD_SIZE 16 
`define ADDR_SIZE 8

//instructions
`define NOP  5'h0
`define LOAD 5'h1
`define STO  5'h2
`define MOV  5'h3
`define ADD  5'h4
`define SUB  5'h5
`define COMP 5'h6
`define JMPU 5'h7
`define JMPC 5'h8
`define MOVG 5'h9
