`define WORD_SIZE 8
