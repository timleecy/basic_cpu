`define WORD_SIZE 8
`define MEM_WIDTH 8 
