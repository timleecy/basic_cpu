`define WORD_SIZE 16 
`define ADDR_SIZE 8

//instructions
`define NOP 5'h0
`define LOADA 5'h1
`define LOADB 5'h2
`define STO 5'h3
